// Computer assembly
//
// Copyright (c) 2025 David Hunter
//
// This program is GPL licensed. See COPYING for the full license.

module mach
  (
   input         CLK,
   input         CE,
   input         RESn,

   output        CPU_BCYSTn,

   output [19:0] ROM_A,
   input [15:0]  ROM_DO,
   output        ROM_CEn,
   input         ROM_READYn,

   output [20:0] RAM_A,
   output [31:0] RAM_DI,
   input [31:0]  RAM_DO,
   output        RAM_CEn,
   output        RAM_WEn,
   output [3:0]  RAM_BEn,
   input         RAM_READYn,

   output [31:0] A
   );

logic [31:0]    dut_ia, dut_da;
logic [31:0]    dut_id;
logic           dut_ireq, dut_iack;
wire [31:0]     dut_dd_i, dut_dd_o;
wire [1:0]      dut_dbc;
wire [3:0]      dut_dbe;
wire            dut_dwr;
wire            dut_dmrq;
wire [1:0]      dut_dst;
wire            dut_dreq, dut_dack;

wire [31:0]     mem_a;
logic [31:0]    mem_d_i;
wire [31:0]     mem_d_o;
wire [3:0]      mem_ben;
wire [1:0]      mem_st;
wire            mem_dan;
wire            mem_mrqn;
wire            mem_rw;
wire            mem_bcystn;
wire            mem_readyn;
wand            mem_szrqn;

logic           rom_cen;
logic [15:0]    rom_do;
logic           rom_readyn;

logic           ram_cen;
wire [31:0]     ram_do;
logic           ram_readyn;

logic           io_cen;
logic           unk_cen;

v810_exec dut
  (
   .RESn(RESn),
   .CLK(CLK),
   .CE(CE),

   .IA(dut_ia),
   .ID(dut_id),
   .IREQ(dut_ireq),
   .IACK(dut_iack),

   .DA(dut_da),
   .DD_I(dut_dd_i),
   .DD_O(dut_dd_o),
   .DBC(dut_dbc),
   .DBE(dut_dbe),
   .DWR(dut_dwr),
   .DMRQ(dut_dmrq),
   .DST(dut_dst),
   .DREQ(dut_dreq),
   .DACK(dut_dack),

   .ST()
   );

v810_mem dut_mem
  (
   .RESn(RESn),
   .CLK(CLK),
   .CE(CE),

   .EUDA(dut_da),
   .EUDD_I(dut_dd_i),
   .EUDD_O(dut_dd_o),
   .EUDBC(dut_dbc),
   .EUDBE(dut_dbe),
   .EUDWR(dut_dwr),
   .EUDMRQ(dut_dmrq),
   .EUDST(dut_dst),
   .EUDREQ(dut_dreq),
   .EUDACK(dut_dack),

   .EUIA(dut_ia),
   .EUID(dut_id),
   .EUIREQ(dut_ireq),
   .EUIACK(dut_iack),

   .A(mem_a),
   .D_I(mem_d_i),
   .D_O(mem_d_o),
   .BEn(mem_ben),
   .ST(mem_st),
   .DAn(mem_dan),
   .MRQn(mem_mrqn),
   .RW(mem_rw),
   .BCYSTn(mem_bcystn),
   .READYn(mem_readyn),
   .SZRQn(mem_szrqn)
   );

always @* begin
    if (~rom_cen)
        mem_d_i = {16'b0, rom_do};
    else if (~ram_cen)
        mem_d_i = ram_do;
    else
        mem_d_i = '0;
end

assign mem_readyn = unk_cen & rom_readyn & ram_readyn & io_cen;
assign mem_szrqn = ~unk_cen | (rom_cen & io_cen);

assign rom_do = ROM_DO;
assign rom_readyn = rom_cen | ROM_READYn;

assign ram_do = RAM_DO;
assign ram_readyn = ram_cen | RAM_READYn;

assign ram_cen = ~(~mem_mrqn & ~mem_a[31]);
assign rom_cen = ~(~mem_mrqn & (mem_a[31:20] == 12'hFFF));
assign io_cen = ~(mem_mrqn & (~mem_bcystn | ~mem_dan) & (mem_st == 2'b10));
assign unk_cen = ~(ram_cen & rom_cen & io_cen);

assign CPU_BCYSTn = mem_bcystn;

assign ROM_CEn = rom_cen;
assign ROM_A = mem_a[19:0];

assign RAM_CEn = ram_cen;
assign RAM_A = mem_a[20:0];
assign RAM_DI = mem_d_o;
assign RAM_WEn = mem_rw;
assign RAM_BEn = mem_ben;

assign A = mem_a;

always @(posedge CLK) if (1 && CE) begin
    if (~io_cen & ~mem_dan)
        $display("%x %s %x", A, (mem_rw ? "R" : "w"),
                 (emem_rw ? mem_d_i[15:0] : mem_d_o[15:0]));
end

endmodule
